----------------------------------------------------------------------------------------------------------------------
-- Title      : Top-level description for <entity>
-- Project    : MUCTPI
----------------------------------------------------------------------------------------------------------------------
-- File       : <filename>
-- Author     : Marcos Oliveira
-- Company    : CERN
-- Created    : <date>
-- Last update: <date>
-- Platform   : Vivado 2016.3 and Mentor Modelsim SE-64 10.1c
-- Standard   : VHDL'93/02
----------------------------------------------------------------------------------------------------------------------
-- Description: Automatically generated with MyPinoutUtils
----------------------------------------------------------------------------------------------------------------------
-- Copyright (c) <year> CERN
----------------------------------------------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- <date>  1.0      msilvaol	Created
----------------------------------------------------------------------------------------------------------------------

entity <entity> is
  port (

end entity <entity>;

architecture rtl of <entity> is

begin  -- architecture rtl

  

end architecture rtl;
