----------------------------------------------------------------------------------------------------------------------
-- Title      : Top-level description for xcvu9pflgc2104pkg
-- Project    : MUCTPI
----------------------------------------------------------------------------------------------------------------------
-- File       : xcvu9pflgc2104pkg_IC15.vhd
-- Author     : Marcos Oliveira
-- Company    : CERN
-- Created    : 2018-11-07
-- Last update: 2018-11-07
-- Platform   : Vivado 2016.3 and Mentor Modelsim SE-64 10.1c
-- Standard   : VHDL'93/02
----------------------------------------------------------------------------------------------------------------------
-- Description: Automatically generated with MyPinoutUtils
----------------------------------------------------------------------------------------------------------------------
-- Copyright (c) 2018 CERN
----------------------------------------------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2018-11-07  1.0      msilvaol	Created
----------------------------------------------------------------------------------------------------------------------

entity xcvu9pflgc2104pkg is
  port (
A2C_DN               : inout std_logic_vector(46 downto 0);
A2C_DP               : inout std_logic_vector(46 downto 0);
C2A_DN               : inout std_logic_vector(46 downto 0);
C2A_DP               : inout std_logic_vector(46 downto 0);
C2T_DN               : inout std_logic_vector(69 downto 0);
C2T_DP               : inout std_logic_vector(69 downto 0);
C2T_GT_N             : inout std_logic_vector(27 downto 0);
C2T_GT_P             : inout std_logic_vector(27 downto 0);
C2Z_AXI_CLK          : inout std_logic;
C2Z_AXI_D            : inout std_logic_vector(21 downto 0);
M2T_MGTCLK_N         : inout std_logic_vector(3 downto 2);
M2T_MGTCLK_P         : inout std_logic_vector(3 downto 2);
MPC_CFG              : inout std_logic_vector(4 downto 0);
MPC_TCK              : inout std_logic;
MPC_TDI              : inout std_logic;
MPC_TMS              : inout std_logic;
SLRX0_N              : inout std_logic_vector(11 downto 0);
SLRX0_P              : inout std_logic_vector(11 downto 0);
SLRX1_N              : inout std_logic_vector(11 downto 0);
SLRX1_P              : inout std_logic_vector(11 downto 0);
SLRX2_N              : inout std_logic_vector(11 downto 0);
SLRX2_P              : inout std_logic_vector(11 downto 0);
SLRX3_N              : inout std_logic_vector(11 downto 0);
SLRX3_P              : inout std_logic_vector(11 downto 0);
SLRX4_N              : inout std_logic_vector(11 downto 0);
SLRX4_P              : inout std_logic_vector(11 downto 0);
SLRX5_N              : inout std_logic_vector(11 downto 0);
SLRX5_P              : inout std_logic_vector(11 downto 0);
SLRX6_N              : inout std_logic_vector(11 downto 0);
SLRX6_P              : inout std_logic_vector(11 downto 0);
SLRX7_N              : inout std_logic_vector(11 downto 0);
SLRX7_P              : inout std_logic_vector(11 downto 0);
SLRX8_N              : inout std_logic_vector(7 downto 0);
SLRX8_P              : inout std_logic_vector(7 downto 0);
SLRX_MGTCLK_N        : inout std_logic_vector(11 downto 6);
SLRX_MGTCLK_P        : inout std_logic_vector(11 downto 6);
SYSMON_AD0_N_C       : inout std_logic;
SYSMON_AD0_P_C       : inout std_logic;
SYSMON_SCL           : inout std_logic_vector(1 downto 1);
SYSMON_SDA           : inout std_logic_vector(1 downto 1);
SYSMON_VN_C          : inout std_logic;
SYSMON_VP_C          : inout std_logic;
SYS_CLK_N            : inout std_logic_vector(1 downto 1);
SYS_CLK_P            : inout std_logic_vector(1 downto 1);
TEMP_DXN_C           : inout std_logic;
TEMP_DXP_C           : inout std_logic;
TPTX0_N              : inout std_logic_vector(11 downto 0);
TPTX0_P              : inout std_logic_vector(11 downto 0);
TPTX1_N              : inout std_logic_vector(11 downto 0);
TPTX1_P              : inout std_logic_vector(11 downto 0);
TPTX_MGTCLK_N        : inout std_logic_vector(3 downto 2);
TPTX_MGTCLK_P        : inout std_logic_vector(3 downto 2);
TP_HPIO71_C          : inout std_logic;
TRP_MPC              : inout std_logic_vector(7 downto 0);
TTC_CLK_N            : inout std_logic_vector(1 downto 1);
TTC_CLK_P            : inout std_logic_vector(1 downto 1);
Z2C_AXI_CLK          : inout std_logic;
Z2C_AXI_D            : inout std_logic_vector(21 downto 0);
ZYQ_CLK_N            : inout std_logic_vector(1 downto 1);
ZYQ_CLK_P            : inout std_logic_vector(1 downto 1);
ZYQ_MPC              : inout std_logic_vector(7 downto 0)
);
end entity xcvu9pflgc2104pkg;

architecture rtl of xcvu9pflgc2104pkg is

begin  -- architecture rtl

  

end architecture rtl;
