----------------------------------------------------------------------------------------------------------------------
-- Title      : Top-level description for <entity>
-- Project    : LASP
----------------------------------------------------------------------------------------------------------------------
-- File       : <filename>
-- Author     : Marcos Oliveira
-- Company    : CERN
-- Created    : <date>
-- Last update: <date>
-- Platform   : Intel Quartus Prime v21.1
-- Standard   : VHDL'93/02
----------------------------------------------------------------------------------------------------------------------
-- Description: Automatically generated with PCBpy
----------------------------------------------------------------------------------------------------------------------
-- Copyright (c) <year> CERN
----------------------------------------------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- <date>  1.0      msilvaol	Created
----------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity <entity> is
  port (

end entity <entity>;

architecture rtl of <entity> is

begin  -- architecture rtl

  

end architecture rtl;
