----------------------------------------------------------------------------------------------------------------------
-- Title      : Top-level description for 1sx280UF50
-- Project    : LASP
----------------------------------------------------------------------------------------------------------------------
-- File       : 1sx280UF50_U4.vhd
-- Author     : Marcos Oliveira
-- Company    : CERN
-- Created    : 2021-04-11
-- Last update: 2021-04-11
-- Platform   : Intel Quartus Prime v21.1
-- Standard   : VHDL'93/02
----------------------------------------------------------------------------------------------------------------------
-- Description: Automatically generated with PCBpy
----------------------------------------------------------------------------------------------------------------------
-- Copyright (c) 2021 CERN
----------------------------------------------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2021-04-11  1.0      msilvaol	Created
----------------------------------------------------------------------------------------------------------------------

entity 1sx280UF50 is
  port (
EXT_STROBE_SX_N      : inout std_logic;
EXT_STROBE_SX_P      : inout std_logic;
FEB_SX_L_N           : inout std_logic_vector(43 downto 0);
FEB_SX_L_P           : inout std_logic_vector(43 downto 0);
FEB_SX_R_N           : inout std_logic_vector(43 downto 0);
FEB_SX_R_P           : inout std_logic_vector(43 downto 0);
FELIX_OPTO_SX_RX_N   : inout std_logic_vector(2 downto 0);
FELIX_OPTO_SX_RX_P   : inout std_logic_vector(2 downto 0);
FELIX_OPTO_SX_TX_N   : inout std_logic_vector(2 downto 0);
FELIX_OPTO_SX_TX_P   : inout std_logic_vector(2 downto 0);
FEX_11_SX_N          : inout std_logic_vector(31 downto 0);
FEX_11_SX_P          : inout std_logic_vector(31 downto 0);
GLOBAL_EV_SX_N       : inout std_logic_vector(3 downto 0);
GLOBAL_EV_SX_P       : inout std_logic_vector(3 downto 0);
HPS_LED01_BLUE_GATE  : inout std_logic;
HPS_LED01_GREEN_GATE : inout std_logic;
HPS_LED01_RED_GATE   : inout std_logic;
HPS_LED02_BLUE_GATE  : inout std_logic;
HPS_LED02_GREEN_GATE : inout std_logic;
HPS_LED02_RED_GATE   : inout std_logic;
HPS_LED03_BLUE_GATE  : inout std_logic;
HPS_LED03_GREEN_GATE : inout std_logic;
HPS_LED03_RED_GATE   : inout std_logic;
HPS_LED04_BLUE_GATE  : inout std_logic;
HPS_LED04_GREEN_GATE : inout std_logic;
HPS_LED04_RED_GATE   : inout std_logic;
HPS_SPI_CLK          : inout std_logic;
HPS_SPI_CS0_N        : inout std_logic;
HPS_SPI_SDO          : inout std_logic;
INPUT_CLK_TO_SX_LEFT_N : inout std_logic;
INPUT_CLK_TO_SX_LEFT_P : inout std_logic;
INPUT_CLK_TO_SX_RIGHT_N : inout std_logic;
INPUT_CLK_TO_SX_RIGHT_P : inout std_logic;
LINK_MAX10_SX_CLK    : inout std_logic;
LINK_MAX10_SX_DATA   : inout std_logic;
LINK_MAX10_SX_VALID  : inout std_logic;
LINK_SX_MAX10_CLK    : inout std_logic;
LINK_SX_MAX10_DATA   : inout std_logic;
LINK_SX_MAX10_VALID  : inout std_logic;
LVDS_CLOCK_TEST_FROM_RTM_SX_AC_N : inout std_logic;
LVDS_CLOCK_TEST_FROM_RTM_SX_AC_P : inout std_logic;
LVDS_CLOCK_TEST_FROM_SX_TO_RTM_N : inout std_logic;
LVDS_CLOCK_TEST_FROM_SX_TO_RTM_P : inout std_logic;
LVDS_DATA_TEST_FROM_RTM_TO_SX_N : inout std_logic;
LVDS_DATA_TEST_FROM_RTM_TO_SX_P : inout std_logic;
LVDS_DATA_TEST_FROM_SX_TO_RTM_N : inout std_logic;
LVDS_DATA_TEST_FROM_SX_TO_RTM_P : inout std_logic;
RCVRD_CLK_FROM_SX_N  : inout std_logic;
RCVRD_CLK_FROM_SX_P  : inout std_logic;
REF_240_SX_LEFT_N    : inout std_logic;
REF_240_SX_LEFT_P    : inout std_logic;
REF_240_SX_RIGHT_N   : inout std_logic;
REF_240_SX_RIGHT_P   : inout std_logic;
RTM_FELIX_SX_AC_RX_N : inout std_logic_vector(0 downto 0);
RTM_FELIX_SX_AC_RX_P : inout std_logic_vector(0 downto 0);
RTM_FELIX_SX_TX_N    : inout std_logic_vector(0 downto 0);
RTM_FELIX_SX_TX_P    : inout std_logic_vector(0 downto 0);
RTM_FEX_25_SX_N      : inout std_logic_vector(19 downto 0);
RTM_FEX_25_SX_P      : inout std_logic_vector(19 downto 0);
RTM_MON_SX_AC_RX_N   : inout std_logic;
RTM_MON_SX_AC_RX_P   : inout std_logic;
RTM_MON_SX_TX_N      : inout std_logic;
RTM_MON_SX_TX_P      : inout std_logic;
SD_CLK               : inout std_logic;
SD_CMD               : inout std_logic;
SD_DATA0             : inout std_logic;
SD_DATA1             : inout std_logic;
SD_DATA2             : inout std_logic;
SD_DATA3             : inout std_logic;
SD_DATA4             : inout std_logic;
SD_DATA5             : inout std_logic;
SD_DATA6             : inout std_logic;
SD_DATA7             : inout std_logic;
SD_PWR_EN            : inout std_logic;
SG210SEH_SX_CLK100_OUT : inout std_logic;
SG210SEH_SX_CLK125_OUT : inout std_logic;
SI530_SX_CLK156_25_N : inout std_logic;
SI530_SX_CLK156_25_P : inout std_logic;
SWITCH_1GBE_SX_RX_N  : inout std_logic;
SWITCH_1GBE_SX_RX_P  : inout std_logic;
SWITCH_1GBE_SX_TX_N  : inout std_logic;
SWITCH_1GBE_SX_TX_P  : inout std_logic;
SX_AS_CLK_R          : inout std_logic;
SX_AS_DATA0          : inout std_logic;
SX_AS_DATA1          : inout std_logic;
SX_AS_DATA2          : inout std_logic;
SX_AS_DATA3          : inout std_logic;
SX_BP0               : inout std_logic;
SX_BP1               : inout std_logic;
SX_CLK_DDR4_COMP_N   : inout std_logic;
SX_CLK_DDR4_COMP_P   : inout std_logic;
SX_CONF_DONE         : inout std_logic;
SX_CONF_INIT_DONE    : inout std_logic;
SX_CONF_NCONFIG      : inout std_logic;
SX_CONF_NSTATUS      : inout std_logic;
SX_CONF_SDM_SCL      : inout std_logic;
SX_CONF_SDM_SDA      : inout std_logic;
SX_DDR4_COMP_A0      : inout std_logic;
SX_DDR4_COMP_A1      : inout std_logic;
SX_DDR4_COMP_A2      : inout std_logic;
SX_DDR4_COMP_A3      : inout std_logic;
SX_DDR4_COMP_A4      : inout std_logic;
SX_DDR4_COMP_A5      : inout std_logic;
SX_DDR4_COMP_A6      : inout std_logic;
SX_DDR4_COMP_A7      : inout std_logic;
SX_DDR4_COMP_A8      : inout std_logic;
SX_DDR4_COMP_A9      : inout std_logic;
SX_DDR4_COMP_A10     : inout std_logic;
SX_DDR4_COMP_A11     : inout std_logic;
SX_DDR4_COMP_A12     : inout std_logic;
SX_DDR4_COMP_A13     : inout std_logic;
SX_DDR4_COMP_A14     : inout std_logic;
SX_DDR4_COMP_A15     : inout std_logic;
SX_DDR4_COMP_A16     : inout std_logic;
SX_DDR4_COMP_ACT_N   : inout std_logic;
SX_DDR4_COMP_ALERT_N : inout std_logic;
SX_DDR4_COMP_BA0     : inout std_logic;
SX_DDR4_COMP_BA1     : inout std_logic;
SX_DDR4_COMP_BG0     : inout std_logic;
SX_DDR4_COMP_BG1     : inout std_logic;
SX_DDR4_COMP_CKE     : inout std_logic;
SX_DDR4_COMP_CLK_N   : inout std_logic;
SX_DDR4_COMP_CLK_P   : inout std_logic;
SX_DDR4_COMP_CS_N    : inout std_logic;
SX_DDR4_COMP_DBI_N0  : inout std_logic;
SX_DDR4_COMP_DBI_N1  : inout std_logic;
SX_DDR4_COMP_DBI_N2  : inout std_logic;
SX_DDR4_COMP_DBI_N3  : inout std_logic;
SX_DDR4_COMP_DQ0     : inout std_logic;
SX_DDR4_COMP_DQ1     : inout std_logic;
SX_DDR4_COMP_DQ2     : inout std_logic;
SX_DDR4_COMP_DQ3     : inout std_logic;
SX_DDR4_COMP_DQ4     : inout std_logic;
SX_DDR4_COMP_DQ5     : inout std_logic;
SX_DDR4_COMP_DQ6     : inout std_logic;
SX_DDR4_COMP_DQ7     : inout std_logic;
SX_DDR4_COMP_DQ8     : inout std_logic;
SX_DDR4_COMP_DQ9     : inout std_logic;
SX_DDR4_COMP_DQ10    : inout std_logic;
SX_DDR4_COMP_DQ11    : inout std_logic;
SX_DDR4_COMP_DQ12    : inout std_logic;
SX_DDR4_COMP_DQ13    : inout std_logic;
SX_DDR4_COMP_DQ14    : inout std_logic;
SX_DDR4_COMP_DQ15    : inout std_logic;
SX_DDR4_COMP_DQ16    : inout std_logic;
SX_DDR4_COMP_DQ17    : inout std_logic;
SX_DDR4_COMP_DQ18    : inout std_logic;
SX_DDR4_COMP_DQ19    : inout std_logic;
SX_DDR4_COMP_DQ20    : inout std_logic;
SX_DDR4_COMP_DQ21    : inout std_logic;
SX_DDR4_COMP_DQ22    : inout std_logic;
SX_DDR4_COMP_DQ23    : inout std_logic;
SX_DDR4_COMP_DQ24    : inout std_logic;
SX_DDR4_COMP_DQ25    : inout std_logic;
SX_DDR4_COMP_DQ26    : inout std_logic;
SX_DDR4_COMP_DQ27    : inout std_logic;
SX_DDR4_COMP_DQ28    : inout std_logic;
SX_DDR4_COMP_DQ29    : inout std_logic;
SX_DDR4_COMP_DQ30    : inout std_logic;
SX_DDR4_COMP_DQ31    : inout std_logic;
SX_DDR4_COMP_DQS_N0  : inout std_logic;
SX_DDR4_COMP_DQS_N1  : inout std_logic;
SX_DDR4_COMP_DQS_N2  : inout std_logic;
SX_DDR4_COMP_DQS_N3  : inout std_logic;
SX_DDR4_COMP_DQS_P0  : inout std_logic;
SX_DDR4_COMP_DQS_P1  : inout std_logic;
SX_DDR4_COMP_DQS_P2  : inout std_logic;
SX_DDR4_COMP_DQS_P3  : inout std_logic;
SX_DDR4_COMP_ODT     : inout std_logic;
SX_DDR4_COMP_PAR     : inout std_logic;
SX_DDR4_COMP_RESET_N : inout std_logic;
SX_DDR4_RZQ          : inout std_logic;
SX_FPGA_TO_RTM_FPGA_GP : inout std_logic;
SX_GP_TEST_IN        : inout std_logic;
SX_GP_TEST_OUT       : inout std_logic;
SX_LED01_BLUE_GATE   : inout std_logic;
SX_LED01_GREEN_GATE  : inout std_logic;
SX_LED01_RED_GATE    : inout std_logic;
SX_LED02_BLUE_GATE   : inout std_logic;
SX_LED02_GREEN_GATE  : inout std_logic;
SX_LED02_RED_GATE    : inout std_logic;
SX_LED03_BLUE_GATE   : inout std_logic;
SX_LED03_GREEN_GATE  : inout std_logic;
SX_LED03_RED_GATE    : inout std_logic;
SX_LED04_BLUE_GATE   : inout std_logic;
SX_LED04_GREEN_GATE  : inout std_logic;
SX_LED04_RED_GATE    : inout std_logic;
SX_LS01_FPGA_OE      : inout std_logic;
SX_LS02_FPGA_OE      : inout std_logic;
SX_LS03_FPGA_OE      : inout std_logic;
SX_LS04_FPGA_OE      : inout std_logic;
SX_LS05_FPGA_OE      : inout std_logic;
SX_LS06_FPGA_OE      : inout std_logic;
SX_LS07_FPGA_OE      : inout std_logic;
SX_LS08_FPGA_OE      : inout std_logic;
SX_LS09_FPGA_OE      : inout std_logic;
SX_LS10_FPGA_OE      : inout std_logic;
SX_LS11_FPGA_OE      : inout std_logic;
SX_LS12_FPGA_OE      : inout std_logic;
SX_MSEL0             : inout std_logic;
SX_MSEL1             : inout std_logic;
SX_MSEL2             : inout std_logic;
SX_PLL_LEMO_OUT_N    : inout std_logic;
SX_PLL_LEMO_OUT_P    : inout std_logic;
SX_REFCLK_641_OUT0_N : inout std_logic;
SX_REFCLK_641_OUT0_P : inout std_logic;
SX_REFCLK_641_OUT1_N : inout std_logic;
SX_REFCLK_641_OUT1_P : inout std_logic;
SX_REFCLK_641_OUT2_N : inout std_logic;
SX_REFCLK_641_OUT2_P : inout std_logic;
SX_REFCLK_641_OUT3_N : inout std_logic;
SX_REFCLK_641_OUT3_P : inout std_logic;
SX_REFCLK_641_OUT4_N : inout std_logic;
SX_REFCLK_641_OUT4_P : inout std_logic;
SX_REFCLK_641_OUT5_N : inout std_logic;
SX_REFCLK_641_OUT5_P : inout std_logic;
SX_REFCLK_641_OUT6_N : inout std_logic;
SX_REFCLK_641_OUT6_P : inout std_logic;
SX_REFCLK_641_OUT7_N : inout std_logic;
SX_REFCLK_641_OUT7_P : inout std_logic;
SX_RESET_N           : inout std_logic;
SX_RX_G1_F01_INTL    : inout std_logic;
SX_RX_G1_F01_PRESENTL : inout std_logic;
SX_RX_G1_F01_RESETL  : inout std_logic;
SX_RX_G1_F01_SELECTL : inout std_logic;
SX_RX_G1_F02_INTL    : inout std_logic;
SX_RX_G1_F02_PRESENTL : inout std_logic;
SX_RX_G1_F02_RESETL  : inout std_logic;
SX_RX_G1_F02_SELECTL : inout std_logic;
SX_RX_G1_F03_INTL    : inout std_logic;
SX_RX_G1_F03_PRESENTL : inout std_logic;
SX_RX_G1_F03_RESETL  : inout std_logic;
SX_RX_G1_F03_SELECTL : inout std_logic;
SX_RX_G1_F04_INTL    : inout std_logic;
SX_RX_G1_F04_PRESENTL : inout std_logic;
SX_RX_G1_F04_RESETL  : inout std_logic;
SX_RX_G1_F04_SELECTL : inout std_logic;
SX_RX_G2_F01_INTL    : inout std_logic;
SX_RX_G2_F01_PRESENTL : inout std_logic;
SX_RX_G2_F01_RESETL  : inout std_logic;
SX_RX_G2_F01_SELECTL : inout std_logic;
SX_RX_G2_F02_INTL    : inout std_logic;
SX_RX_G2_F02_PRESENTL : inout std_logic;
SX_RX_G2_F02_RESETL  : inout std_logic;
SX_RX_G2_F02_SELECTL : inout std_logic;
SX_RX_G2_F03_INTL    : inout std_logic;
SX_RX_G2_F03_PRESENTL : inout std_logic;
SX_RX_G2_F03_RESETL  : inout std_logic;
SX_RX_G2_F03_SELECTL : inout std_logic;
SX_RX_G2_F04_INTL    : inout std_logic;
SX_RX_G2_F04_PRESENTL : inout std_logic;
SX_RX_G2_F04_RESETL  : inout std_logic;
SX_RX_G2_F04_SELECTL : inout std_logic;
SX_RX_G2_SCL         : inout std_logic;
SX_RX_G2_SDA         : inout std_logic;
SX_TEMPDIODE0_N      : inout std_logic;
SX_TEMPDIODE0_P      : inout std_logic;
SX_TEMPDIODE1_N      : inout std_logic;
SX_TEMPDIODE1_P      : inout std_logic;
SX_TEST_CLK_IN0_N    : inout std_logic;
SX_TEST_CLK_IN0_P    : inout std_logic;
SX_TEST_CLK_IN1_N    : inout std_logic;
SX_TEST_CLK_IN1_P    : inout std_logic;
SX_TEST_CLK_OUT0_N   : inout std_logic;
SX_TEST_CLK_OUT0_P   : inout std_logic;
SX_TEST_CLK_OUT1_N   : inout std_logic;
SX_TEST_CLK_OUT1_P   : inout std_logic;
SX_TX_G1_F01_INTL    : inout std_logic;
SX_TX_G1_F01_PRESENTL : inout std_logic;
SX_TX_G1_F01_RESETL  : inout std_logic;
SX_TX_G1_F01_SELECTL : inout std_logic;
SX_TX_G1_F02_INTL    : inout std_logic;
SX_TX_G1_F02_PRESENTL : inout std_logic;
SX_TX_G1_F02_RESETL  : inout std_logic;
SX_TX_G1_F02_SELECTL : inout std_logic;
SX_TX_G1_F03_INTL    : inout std_logic;
SX_TX_G1_F03_PRESENTL : inout std_logic;
SX_TX_G1_F03_RESETL  : inout std_logic;
SX_TX_G1_F03_SELECTL : inout std_logic;
SX_TX_G1_F04_INTL    : inout std_logic;
SX_TX_G1_F04_PRESENTL : inout std_logic;
SX_TX_G1_F04_RESETL  : inout std_logic;
SX_TX_G1_F04_SELECTL : inout std_logic;
SX_TX_RX_G1_SCL      : inout std_logic;
SX_TX_RX_G1_SDA      : inout std_logic;
SX_USER0             : inout std_logic;
SX_USER1             : inout std_logic;
SX_USER2             : inout std_logic;
SX_USER3             : inout std_logic;
SX_VCXO_DOWN         : inout std_logic;
SX_VCXO_UP           : inout std_logic;
TCK_FOR_SX           : inout std_logic;
TDI_FOR_SX           : inout std_logic;
TDO_FOR_SX           : inout std_logic;
TMS_FOR_SX           : inout std_logic
);
end entity 1sx280UF50;

architecture rtl of 1sx280UF50 is

begin  -- architecture rtl

  

end architecture rtl;
